module sq_wave_gen (
    input clk,
    input next_sample,
    output [9:0] code
);

    // Remove this line once you create your square wave generator
    assign code = 0;
endmodule

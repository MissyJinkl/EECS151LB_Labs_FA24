module nco(
    input clk,
    input rst,
    input [23:0] fcw,
    input next_sample,
    output [9:0] code
);

    // Remove this line once you create your nco
    assign code = 0;
endmodule
